library ieee;
use ieee.std_logic_1164.all;
use work.definitions.all;

entity fib_generator is
-- 	port (
-- 		out_fwd : in channel_forward;
-- 		out_bck : out channel_backward	
-- 	);
end entity fib_generator;


architecture struct of fib_generator is
begin
	
	-- TODO

end architecture struct;

